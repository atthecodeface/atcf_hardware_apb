/** Copyright (C) 2016-2017,  Gavin J Stark.  All rights reserved.
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *   http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * @file  tb_apb_processor.cdl
 * @brief Testbench for APB processor (ROM-based APB trasanctions)
 *
 * This is a simple testbench for the ROM-based APB transaction processor
 */
/*a Includes */
include "std::srams.h"
include "apb.h"
include "apb_utilities.h"
include "apb_targets.h"
include "apb_masters.h"

/*a Module */
module tb_apb_processor( clock clk,
                         input bit reset_n,
                         input t_apb_processor_request  apb_processor_request,
                         output t_apb_processor_response  apb_processor_response,
                         output bit[3] timer_equalled
)
{

    /*b Nets */
    net t_apb_processor_response  apb_processor_response;
    net t_apb_request             apb_request;
    net t_apb_rom_request         rom_request;
    net bit[40]                   rom_data;
    net t_apb_response timer_apb_response;
    net t_apb_response gpio_apb_response;
    net bit[3] timer_equalled;
    comb t_apb_response            apb_response;
    comb t_apb_request timer_apb_request;
    comb t_apb_request gpio_apb_request;

    net bit[16] gpio_output;
    net bit[16] gpio_output_enable;
    comb bit[16]  gpio_input;
    net bit     gpio_input_event;

    /*b Instantiations */
    instantiations: {
        apb_processor apbp( clk <- clk,
                       reset_n <= reset_n,

                       apb_processor_request <= apb_processor_request,
                       apb_processor_response => apb_processor_response,
                       apb_request => apb_request,
                       apb_response  <= apb_response,
                       rom_request => rom_request,
                       rom_data <= rom_data );

        se_sram_srw_16384x40 apb_rom(sram_clock <- clk,
                                     select <= rom_request.enable,
                                     address <= rom_request.address[14;0],
                                     read_not_write <= 1,
                                     write_data <= 0,
                                     data_out => rom_data );

        apb_target_timer timer( clk <- clk,
                                reset_n <= reset_n,
                                apb_request  <= timer_apb_request,
                                apb_response => timer_apb_response,
                                timer_equalled => timer_equalled );

        apb_target_gpio gpio( clk <- clk,
                              reset_n <= reset_n,
                              apb_request  <= gpio_apb_request,
                              apb_response => gpio_apb_response,
                              gpio_input <= gpio_input,
                              gpio_output => gpio_output,
                              gpio_output_enable => gpio_output_enable,
                              gpio_input_event => gpio_input_event
            );
        timer_apb_request = apb_request;
        gpio_apb_request = apb_request;
        timer_apb_request.psel = apb_request.psel && (apb_request.paddr[4;28]==0);
        gpio_apb_request.psel  = apb_request.psel && (apb_request.paddr[4;28]==1);
        apb_response = timer_apb_response;
        if (apb_request.paddr[4;28]==1) { apb_response = gpio_apb_response; }
        gpio_input = bundle(13b0, timer_equalled);
    }

    /*b Logging */
    default clock clk;
    default reset active_low reset_n;
    clocked t_apb_rom_request log_rom_request={*=0};
    logging : {
        apb_logging apb_log( clk <- clk, reset_n <= reset_n, apb_request <= apb_request, apb_response <= apb_response );
        log_rom_request <= rom_request;
        if (log_rom_request.enable) {
            log("sram_read", "address", log_rom_request.address, "data", rom_data );
        }
    }

    /*b All done */
}
